module and_gate (input a, input b, output y);//data flow mmodelling 
  assign y = a & b;
endmodule
